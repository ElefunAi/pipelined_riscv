module sample_test ();
// build/c_sample.hex
    
endmodule